`timescale 1ns/10ps
module immediate_offset_unit (
);

endmodule
